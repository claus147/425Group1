----------------------------------------------------------------------------------------
-- This module is used hold values inbetween EX_MEM (Buffer)
-- 
-- Inputs:
-- - ALUE, ALU output
-- - RdtE, register name (for forwarding)
-- - MemReadE
-- - MemWriteE
-- - MemtoRegE
-- - RegWriteE
-- - DumpE, Main_Memory line
-- - ResetE, Main_Memory line
-- - InitMemE, Main_Memory line
-- - WordByteE, Main_Memory line
--
-- Outputs:						
-- - ALUW, ALU output
-- - RdtW, register name (for forwarding)
-- - MemReadW
-- - MemWriteW
-- - MemtoRegW
-- - RegWriteW
-- - DumpW, Main_Memory line
-- - ResetW, Main_Memory line
-- - InitMemW, Main_Memory line
-- - WordByteW, Main_Memory line
--	
-- Control:
-- 	- clk		clock
-- 
--
----------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
----------------------------------------------------------------
entity Reg_EX_MEM is
	port (
		clk 				: in std_logic;
		rst 				: in std_logic;
		ALUE    : in signed(31 downto 0);
		ALUM    : out signed(31 downto 0);
	  RdtE    : in std_ulogic_vector(4 downto 0);
		RdtM    : out std_ulogic_vector(4 downto 0);
    MemWriteE, MemtoRegE,RegWriteE,WordByteE : in std_logic;
	  MemWriteM, MemtoRegM,RegWriteM,WordByteM : out std_logic;
	  WriteDataE : in signed(31 downto 0);
	  writeDataM	: out  signed(31 downto 0)
	);
end entity Reg_EX_MEM;
--------------------------------------------------------------
architecture RTL of Reg_EX_MEM is
  
begin
  process(clk,rst)
  begin
   if (rst = '1') then
 	  ALUM <= (OTHERS => '0');
	  MemWriteM <= '0';
	  MemtoRegM <= '0';
	  RegWriteM <= '0';
	  WordByteM <= '1';
	  RdtM <= (OTHERS => '0');
	  WriteDataM <= (OTHERS => '0');
	 elsif(rising_edge(clk)) then 
	  ALUM <= ALUE;
	  MemWriteM <= MemWriteE;
	  MemtoRegM <= MemtoRegE; 
	  RegWriteM <= RegWriteE;
	  WordByteM <= WordByteE;
	  RdtM <= RdtE;
	  WriteDataM <= WriteDataE;
	 end if;
	end process;   

end architecture RTL;


